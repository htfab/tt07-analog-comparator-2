VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Saitama224_comp
  CLASS BLOCK ;
  FOREIGN tt_um_Saitama224_comp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.600000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 9.816400 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 137.740 11.465 139.850 14.655 ;
        RECT 142.790 11.435 154.060 14.625 ;
      LAYER pwell ;
        RECT 137.670 7.165 139.780 10.265 ;
        RECT 142.690 8.065 153.960 10.300 ;
        RECT 142.430 7.825 153.960 8.065 ;
        RECT 142.690 7.200 153.960 7.825 ;
      LAYER li1 ;
        RECT 138.460 14.475 139.135 14.520 ;
        RECT 137.920 14.305 139.670 14.475 ;
        RECT 143.825 14.445 152.985 14.595 ;
        RECT 137.920 11.815 138.090 14.305 ;
        RECT 138.460 14.245 139.135 14.305 ;
        RECT 138.630 13.795 138.960 13.965 ;
        RECT 138.490 12.540 138.660 13.580 ;
        RECT 138.930 12.540 139.100 13.580 ;
        RECT 138.630 12.155 138.960 12.325 ;
        RECT 139.500 11.815 139.670 14.305 ;
        RECT 137.920 11.645 139.670 11.815 ;
        RECT 142.970 14.275 153.880 14.445 ;
        RECT 142.970 11.785 143.140 14.275 ;
        RECT 143.825 14.245 152.985 14.275 ;
        RECT 144.180 13.765 144.510 13.935 ;
        RECT 145.140 13.765 145.470 13.935 ;
        RECT 146.100 13.765 146.430 13.935 ;
        RECT 147.060 13.765 147.390 13.935 ;
        RECT 148.020 13.765 148.350 13.935 ;
        RECT 148.980 13.765 149.310 13.935 ;
        RECT 149.940 13.765 150.270 13.935 ;
        RECT 150.900 13.765 151.230 13.935 ;
        RECT 151.860 13.765 152.190 13.935 ;
        RECT 152.820 13.765 153.150 13.935 ;
        RECT 143.540 12.510 143.710 13.550 ;
        RECT 144.020 12.510 144.190 13.550 ;
        RECT 144.500 12.510 144.670 13.550 ;
        RECT 144.980 12.510 145.150 13.550 ;
        RECT 145.460 12.510 145.630 13.550 ;
        RECT 145.940 12.510 146.110 13.550 ;
        RECT 146.420 12.510 146.590 13.550 ;
        RECT 146.900 12.510 147.070 13.550 ;
        RECT 147.380 12.510 147.550 13.550 ;
        RECT 147.860 12.510 148.030 13.550 ;
        RECT 148.340 12.510 148.510 13.550 ;
        RECT 148.820 12.510 148.990 13.550 ;
        RECT 149.300 12.510 149.470 13.550 ;
        RECT 149.780 12.510 149.950 13.550 ;
        RECT 150.260 12.510 150.430 13.550 ;
        RECT 150.740 12.510 150.910 13.550 ;
        RECT 151.220 12.510 151.390 13.550 ;
        RECT 151.700 12.510 151.870 13.550 ;
        RECT 152.180 12.510 152.350 13.550 ;
        RECT 152.660 12.510 152.830 13.550 ;
        RECT 153.140 12.510 153.310 13.550 ;
        RECT 143.700 12.125 144.030 12.295 ;
        RECT 144.660 12.125 144.990 12.295 ;
        RECT 145.620 12.125 145.950 12.295 ;
        RECT 146.580 12.125 146.910 12.295 ;
        RECT 147.540 12.125 147.870 12.295 ;
        RECT 148.500 12.125 148.830 12.295 ;
        RECT 149.460 12.125 149.790 12.295 ;
        RECT 150.420 12.125 150.750 12.295 ;
        RECT 151.380 12.125 151.710 12.295 ;
        RECT 152.340 12.125 152.670 12.295 ;
        RECT 153.710 11.785 153.880 14.275 ;
        RECT 142.970 11.615 153.880 11.785 ;
        RECT 137.850 9.915 139.600 10.085 ;
        RECT 137.850 7.515 138.020 9.915 ;
        RECT 138.560 9.405 138.890 9.575 ;
        RECT 138.420 8.195 138.590 9.235 ;
        RECT 138.860 8.195 139.030 9.235 ;
        RECT 138.560 7.855 138.890 8.025 ;
        RECT 138.405 7.515 139.080 7.580 ;
        RECT 139.430 7.515 139.600 9.915 ;
        RECT 137.850 7.345 139.600 7.515 ;
        RECT 142.870 9.950 153.780 10.120 ;
        RECT 142.870 7.550 143.040 9.950 ;
        RECT 144.080 9.440 144.410 9.610 ;
        RECT 145.040 9.440 145.370 9.610 ;
        RECT 146.000 9.440 146.330 9.610 ;
        RECT 146.960 9.440 147.290 9.610 ;
        RECT 147.920 9.440 148.250 9.610 ;
        RECT 148.880 9.440 149.210 9.610 ;
        RECT 149.840 9.440 150.170 9.610 ;
        RECT 150.800 9.440 151.130 9.610 ;
        RECT 151.760 9.440 152.090 9.610 ;
        RECT 152.720 9.440 153.050 9.610 ;
        RECT 143.440 8.230 143.610 9.270 ;
        RECT 143.920 8.230 144.090 9.270 ;
        RECT 144.400 8.230 144.570 9.270 ;
        RECT 144.880 8.230 145.050 9.270 ;
        RECT 145.360 8.230 145.530 9.270 ;
        RECT 145.840 8.230 146.010 9.270 ;
        RECT 146.320 8.230 146.490 9.270 ;
        RECT 146.800 8.230 146.970 9.270 ;
        RECT 147.280 8.230 147.450 9.270 ;
        RECT 147.760 8.230 147.930 9.270 ;
        RECT 148.240 8.230 148.410 9.270 ;
        RECT 148.720 8.230 148.890 9.270 ;
        RECT 149.200 8.230 149.370 9.270 ;
        RECT 149.680 8.230 149.850 9.270 ;
        RECT 150.160 8.230 150.330 9.270 ;
        RECT 150.640 8.230 150.810 9.270 ;
        RECT 151.120 8.230 151.290 9.270 ;
        RECT 151.600 8.230 151.770 9.270 ;
        RECT 152.080 8.230 152.250 9.270 ;
        RECT 152.560 8.230 152.730 9.270 ;
        RECT 153.040 8.230 153.210 9.270 ;
        RECT 143.600 7.890 143.930 8.060 ;
        RECT 144.560 7.890 144.890 8.060 ;
        RECT 145.520 7.890 145.850 8.060 ;
        RECT 146.480 7.890 146.810 8.060 ;
        RECT 147.440 7.890 147.770 8.060 ;
        RECT 148.400 7.890 148.730 8.060 ;
        RECT 149.360 7.890 149.690 8.060 ;
        RECT 150.320 7.890 150.650 8.060 ;
        RECT 151.280 7.890 151.610 8.060 ;
        RECT 152.240 7.890 152.570 8.060 ;
        RECT 143.840 7.550 153.000 7.605 ;
        RECT 153.610 7.550 153.780 9.950 ;
        RECT 142.870 7.380 153.780 7.550 ;
        RECT 138.405 7.305 139.080 7.345 ;
        RECT 143.840 7.255 153.000 7.380 ;
      LAYER met1 ;
        RECT 129.700 16.960 131.200 16.990 ;
        RECT 129.700 16.550 135.990 16.960 ;
        RECT 129.700 15.550 156.660 16.550 ;
        RECT 129.700 15.460 136.745 15.550 ;
        RECT 129.700 15.430 131.200 15.460 ;
        RECT 135.975 12.665 136.745 15.460 ;
        RECT 138.295 14.160 139.295 15.550 ;
        RECT 137.095 13.985 137.315 14.000 ;
        RECT 138.650 13.985 138.940 13.995 ;
        RECT 137.095 13.765 138.980 13.985 ;
        RECT 137.095 12.350 137.315 13.765 ;
        RECT 141.580 13.595 141.920 15.550 ;
        RECT 143.645 14.175 153.155 15.550 ;
        RECT 142.400 13.725 153.210 13.965 ;
        RECT 138.460 13.465 138.690 13.560 ;
        RECT 138.900 13.475 139.130 13.560 ;
        RECT 137.660 12.695 138.700 13.465 ;
        RECT 138.460 12.560 138.690 12.695 ;
        RECT 138.870 12.665 140.775 13.475 ;
        RECT 141.550 13.255 141.950 13.595 ;
        RECT 138.900 12.560 139.130 12.665 ;
        RECT 138.650 12.350 138.940 12.355 ;
        RECT 137.095 12.130 138.970 12.350 ;
        RECT 134.330 11.280 135.230 11.290 ;
        RECT 134.330 10.885 136.070 11.280 ;
        RECT 137.095 10.885 137.315 12.130 ;
        RECT 138.650 12.125 138.940 12.130 ;
        RECT 134.330 10.665 137.315 10.885 ;
        RECT 134.330 10.340 136.070 10.665 ;
        RECT 134.300 10.280 136.070 10.340 ;
        RECT 134.300 9.440 135.260 10.280 ;
        RECT 137.095 9.590 137.315 10.665 ;
        RECT 139.965 11.180 140.775 12.665 ;
        RECT 142.400 12.305 142.640 13.725 ;
        RECT 143.420 13.285 143.820 13.575 ;
        RECT 143.510 12.530 143.740 13.285 ;
        RECT 143.990 12.855 144.220 13.530 ;
        RECT 144.390 13.275 144.790 13.565 ;
        RECT 143.900 12.565 144.300 12.855 ;
        RECT 143.990 12.530 144.220 12.565 ;
        RECT 144.470 12.530 144.700 13.275 ;
        RECT 144.950 12.865 145.180 13.530 ;
        RECT 145.360 13.275 145.760 13.565 ;
        RECT 144.860 12.575 145.260 12.865 ;
        RECT 144.950 12.530 145.180 12.575 ;
        RECT 145.430 12.530 145.660 13.275 ;
        RECT 145.910 12.855 146.140 13.530 ;
        RECT 146.310 13.275 146.710 13.565 ;
        RECT 145.820 12.565 146.220 12.855 ;
        RECT 145.910 12.530 146.140 12.565 ;
        RECT 146.390 12.530 146.620 13.275 ;
        RECT 146.870 12.855 147.100 13.530 ;
        RECT 147.260 13.275 147.660 13.565 ;
        RECT 146.780 12.565 147.180 12.855 ;
        RECT 146.870 12.530 147.100 12.565 ;
        RECT 147.350 12.530 147.580 13.275 ;
        RECT 147.830 12.855 148.060 13.530 ;
        RECT 148.220 13.275 148.620 13.565 ;
        RECT 147.740 12.565 148.140 12.855 ;
        RECT 147.830 12.530 148.060 12.565 ;
        RECT 148.310 12.530 148.540 13.275 ;
        RECT 148.790 12.865 149.020 13.530 ;
        RECT 149.190 13.285 149.590 13.575 ;
        RECT 148.690 12.575 149.090 12.865 ;
        RECT 148.790 12.530 149.020 12.575 ;
        RECT 149.270 12.530 149.500 13.285 ;
        RECT 149.750 12.855 149.980 13.530 ;
        RECT 150.140 13.275 150.540 13.565 ;
        RECT 149.660 12.565 150.060 12.855 ;
        RECT 149.750 12.530 149.980 12.565 ;
        RECT 150.230 12.530 150.460 13.275 ;
        RECT 150.710 12.855 150.940 13.530 ;
        RECT 151.110 13.285 151.510 13.575 ;
        RECT 150.620 12.565 151.020 12.855 ;
        RECT 150.710 12.530 150.940 12.565 ;
        RECT 151.190 12.530 151.420 13.285 ;
        RECT 151.670 12.855 151.900 13.530 ;
        RECT 152.060 13.285 152.460 13.575 ;
        RECT 151.570 12.565 151.970 12.855 ;
        RECT 151.670 12.530 151.900 12.565 ;
        RECT 152.150 12.530 152.380 13.285 ;
        RECT 152.630 12.855 152.860 13.530 ;
        RECT 153.030 13.275 153.430 13.565 ;
        RECT 152.540 12.565 152.940 12.855 ;
        RECT 152.630 12.530 152.860 12.565 ;
        RECT 153.110 12.530 153.340 13.275 ;
        RECT 154.380 12.555 154.780 12.895 ;
        RECT 143.720 12.305 144.010 12.325 ;
        RECT 144.680 12.305 144.970 12.325 ;
        RECT 145.640 12.305 145.930 12.325 ;
        RECT 146.600 12.305 146.890 12.325 ;
        RECT 147.560 12.305 147.850 12.325 ;
        RECT 148.520 12.305 148.810 12.325 ;
        RECT 149.480 12.305 149.770 12.325 ;
        RECT 150.440 12.305 150.730 12.325 ;
        RECT 151.400 12.305 151.690 12.325 ;
        RECT 152.360 12.305 152.650 12.325 ;
        RECT 142.400 12.065 153.230 12.305 ;
        RECT 142.400 11.180 142.640 12.065 ;
        RECT 139.965 10.370 142.640 11.180 ;
        RECT 154.410 10.955 154.750 12.555 ;
        RECT 156.410 11.280 157.310 11.330 ;
        RECT 155.655 10.955 157.310 11.280 ;
        RECT 154.410 10.875 157.310 10.955 ;
        RECT 138.580 9.590 138.870 9.605 ;
        RECT 137.095 9.370 138.905 9.590 ;
        RECT 129.690 6.610 131.190 6.640 ;
        RECT 129.690 6.400 135.660 6.610 ;
        RECT 135.955 6.400 136.745 9.125 ;
        RECT 137.095 8.050 137.315 9.370 ;
        RECT 138.390 9.095 138.620 9.215 ;
        RECT 138.830 9.110 139.060 9.215 ;
        RECT 139.965 9.110 140.775 10.370 ;
        RECT 137.590 8.305 138.630 9.095 ;
        RECT 138.390 8.215 138.620 8.305 ;
        RECT 138.825 8.300 140.775 9.110 ;
        RECT 142.400 9.635 142.640 10.370 ;
        RECT 154.380 10.615 157.310 10.875 ;
        RECT 154.380 10.605 154.750 10.615 ;
        RECT 144.100 9.635 144.390 9.640 ;
        RECT 145.060 9.635 145.350 9.640 ;
        RECT 146.020 9.635 146.310 9.640 ;
        RECT 146.980 9.635 147.270 9.640 ;
        RECT 147.940 9.635 148.230 9.640 ;
        RECT 148.900 9.635 149.190 9.640 ;
        RECT 149.860 9.635 150.150 9.640 ;
        RECT 150.820 9.635 151.110 9.640 ;
        RECT 151.780 9.635 152.070 9.640 ;
        RECT 152.740 9.635 153.030 9.640 ;
        RECT 142.400 9.395 153.240 9.635 ;
        RECT 138.830 8.215 139.060 8.300 ;
        RECT 141.550 8.265 141.950 8.605 ;
        RECT 138.580 8.050 138.870 8.055 ;
        RECT 137.095 7.830 138.870 8.050 ;
        RECT 138.580 7.825 138.870 7.830 ;
        RECT 138.235 6.400 139.235 7.645 ;
        RECT 141.580 6.400 141.920 8.265 ;
        RECT 142.400 8.065 142.640 9.395 ;
        RECT 154.380 9.275 154.720 10.605 ;
        RECT 155.655 10.370 157.310 10.615 ;
        RECT 155.655 10.280 157.340 10.370 ;
        RECT 156.380 9.470 157.340 10.280 ;
        RECT 143.410 8.575 143.640 9.250 ;
        RECT 143.890 9.245 144.120 9.250 ;
        RECT 143.810 8.955 144.210 9.245 ;
        RECT 143.320 8.285 143.720 8.575 ;
        RECT 143.410 8.250 143.640 8.285 ;
        RECT 143.890 8.250 144.120 8.955 ;
        RECT 144.370 8.575 144.600 9.250 ;
        RECT 144.850 9.245 145.080 9.250 ;
        RECT 144.760 8.955 145.160 9.245 ;
        RECT 144.280 8.285 144.680 8.575 ;
        RECT 144.370 8.250 144.600 8.285 ;
        RECT 144.850 8.250 145.080 8.955 ;
        RECT 145.330 8.575 145.560 9.250 ;
        RECT 145.810 9.245 146.040 9.250 ;
        RECT 145.730 8.955 146.130 9.245 ;
        RECT 145.250 8.285 145.650 8.575 ;
        RECT 145.330 8.250 145.560 8.285 ;
        RECT 145.810 8.250 146.040 8.955 ;
        RECT 146.290 8.565 146.520 9.250 ;
        RECT 146.680 8.965 147.080 9.255 ;
        RECT 146.200 8.275 146.600 8.565 ;
        RECT 146.290 8.250 146.520 8.275 ;
        RECT 146.770 8.250 147.000 8.965 ;
        RECT 147.250 8.575 147.480 9.250 ;
        RECT 147.650 8.965 148.050 9.255 ;
        RECT 147.170 8.285 147.570 8.575 ;
        RECT 147.250 8.250 147.480 8.285 ;
        RECT 147.730 8.250 147.960 8.965 ;
        RECT 148.210 8.575 148.440 9.250 ;
        RECT 148.610 8.965 149.010 9.255 ;
        RECT 148.120 8.285 148.520 8.575 ;
        RECT 148.210 8.250 148.440 8.285 ;
        RECT 148.690 8.250 148.920 8.965 ;
        RECT 149.170 8.575 149.400 9.250 ;
        RECT 149.650 9.245 149.880 9.250 ;
        RECT 149.570 8.955 149.970 9.245 ;
        RECT 149.080 8.285 149.480 8.575 ;
        RECT 149.170 8.250 149.400 8.285 ;
        RECT 149.650 8.250 149.880 8.955 ;
        RECT 150.130 8.575 150.360 9.250 ;
        RECT 150.610 9.245 150.840 9.250 ;
        RECT 150.530 8.955 150.930 9.245 ;
        RECT 150.050 8.285 150.450 8.575 ;
        RECT 150.130 8.250 150.360 8.285 ;
        RECT 150.610 8.250 150.840 8.955 ;
        RECT 151.090 8.575 151.320 9.250 ;
        RECT 151.570 9.245 151.800 9.250 ;
        RECT 151.490 8.955 151.890 9.245 ;
        RECT 151.000 8.285 151.400 8.575 ;
        RECT 151.090 8.250 151.320 8.285 ;
        RECT 151.570 8.250 151.800 8.955 ;
        RECT 152.050 8.585 152.280 9.250 ;
        RECT 152.530 9.235 152.760 9.250 ;
        RECT 152.450 8.945 152.850 9.235 ;
        RECT 151.980 8.295 152.380 8.585 ;
        RECT 152.050 8.250 152.280 8.295 ;
        RECT 152.530 8.250 152.760 8.945 ;
        RECT 153.010 8.575 153.240 9.250 ;
        RECT 154.350 8.935 154.750 9.275 ;
        RECT 152.930 8.285 153.330 8.575 ;
        RECT 153.010 8.250 153.240 8.285 ;
        RECT 143.620 8.065 143.910 8.090 ;
        RECT 144.580 8.065 144.870 8.090 ;
        RECT 145.540 8.065 145.830 8.090 ;
        RECT 146.500 8.065 146.790 8.090 ;
        RECT 147.460 8.065 147.750 8.090 ;
        RECT 148.420 8.065 148.710 8.090 ;
        RECT 149.380 8.065 149.670 8.090 ;
        RECT 150.340 8.065 150.630 8.090 ;
        RECT 151.300 8.065 151.590 8.090 ;
        RECT 152.260 8.065 152.550 8.090 ;
        RECT 142.400 7.825 153.240 8.065 ;
        RECT 143.575 6.400 153.210 7.675 ;
        RECT 129.690 5.400 156.630 6.400 ;
        RECT 129.690 5.110 135.660 5.400 ;
        RECT 129.690 5.080 131.190 5.110 ;
      LAYER met2 ;
        RECT 126.735 16.960 128.185 16.980 ;
        RECT 126.710 15.460 131.230 16.960 ;
        RECT 126.735 15.440 128.185 15.460 ;
        RECT 141.580 13.595 141.920 13.625 ;
        RECT 143.470 13.595 143.770 13.625 ;
        RECT 144.440 13.595 144.740 13.615 ;
        RECT 145.410 13.595 145.710 13.615 ;
        RECT 146.360 13.595 146.660 13.615 ;
        RECT 147.310 13.595 147.610 13.615 ;
        RECT 148.270 13.595 148.570 13.615 ;
        RECT 149.240 13.595 149.540 13.625 ;
        RECT 150.190 13.595 150.490 13.615 ;
        RECT 151.160 13.595 151.460 13.625 ;
        RECT 152.110 13.595 152.410 13.625 ;
        RECT 153.080 13.595 153.380 13.615 ;
        RECT 137.690 13.465 138.460 13.495 ;
        RECT 135.945 12.695 138.460 13.465 ;
        RECT 141.580 13.255 153.540 13.595 ;
        RECT 141.580 13.225 141.920 13.255 ;
        RECT 143.470 13.235 143.770 13.255 ;
        RECT 144.440 13.225 144.740 13.255 ;
        RECT 145.410 13.225 145.710 13.255 ;
        RECT 146.360 13.225 146.660 13.255 ;
        RECT 147.310 13.225 147.610 13.255 ;
        RECT 148.270 13.225 148.570 13.255 ;
        RECT 149.240 13.235 149.540 13.255 ;
        RECT 150.190 13.225 150.490 13.255 ;
        RECT 151.160 13.235 151.460 13.255 ;
        RECT 152.110 13.235 152.410 13.255 ;
        RECT 153.080 13.225 153.380 13.255 ;
        RECT 143.950 12.895 144.250 12.905 ;
        RECT 144.910 12.895 145.210 12.915 ;
        RECT 145.870 12.895 146.170 12.905 ;
        RECT 146.830 12.895 147.130 12.905 ;
        RECT 147.790 12.895 148.090 12.905 ;
        RECT 148.740 12.895 149.040 12.915 ;
        RECT 149.710 12.895 150.010 12.905 ;
        RECT 150.670 12.895 150.970 12.905 ;
        RECT 151.620 12.895 151.920 12.905 ;
        RECT 152.590 12.895 152.890 12.905 ;
        RECT 154.410 12.895 154.750 12.925 ;
        RECT 137.690 12.665 138.460 12.695 ;
        RECT 141.570 12.555 154.750 12.895 ;
        RECT 143.950 12.515 144.250 12.555 ;
        RECT 144.910 12.525 145.210 12.555 ;
        RECT 145.870 12.515 146.170 12.555 ;
        RECT 146.830 12.515 147.130 12.555 ;
        RECT 147.790 12.515 148.090 12.555 ;
        RECT 148.740 12.525 149.040 12.555 ;
        RECT 149.710 12.515 150.010 12.555 ;
        RECT 150.670 12.515 150.970 12.555 ;
        RECT 151.620 12.515 151.920 12.555 ;
        RECT 152.590 12.515 152.890 12.555 ;
        RECT 154.410 12.525 154.750 12.555 ;
        RECT 134.330 9.395 135.230 10.370 ;
        RECT 134.310 8.545 135.250 9.395 ;
        RECT 156.410 9.365 157.310 10.400 ;
        RECT 143.860 9.275 144.160 9.295 ;
        RECT 144.810 9.275 145.110 9.295 ;
        RECT 145.780 9.275 146.080 9.295 ;
        RECT 146.730 9.275 147.030 9.305 ;
        RECT 147.700 9.275 148.000 9.305 ;
        RECT 148.660 9.275 148.960 9.305 ;
        RECT 149.620 9.275 149.920 9.295 ;
        RECT 150.580 9.275 150.880 9.295 ;
        RECT 151.540 9.275 151.840 9.295 ;
        RECT 152.500 9.275 152.800 9.285 ;
        RECT 154.380 9.275 154.720 9.305 ;
        RECT 137.620 9.095 138.410 9.125 ;
        RECT 134.330 8.520 135.230 8.545 ;
        RECT 135.925 8.305 138.410 9.095 ;
        RECT 141.580 8.935 154.720 9.275 ;
        RECT 143.860 8.905 144.160 8.935 ;
        RECT 144.810 8.905 145.110 8.935 ;
        RECT 145.780 8.905 146.080 8.935 ;
        RECT 146.730 8.915 147.030 8.935 ;
        RECT 147.700 8.915 148.000 8.935 ;
        RECT 148.660 8.915 148.960 8.935 ;
        RECT 149.620 8.905 149.920 8.935 ;
        RECT 150.580 8.905 150.880 8.935 ;
        RECT 151.540 8.905 151.840 8.935 ;
        RECT 152.500 8.895 152.800 8.935 ;
        RECT 154.380 8.905 154.720 8.935 ;
        RECT 137.620 8.275 138.410 8.305 ;
        RECT 141.580 8.605 141.920 8.635 ;
        RECT 143.370 8.605 143.670 8.625 ;
        RECT 144.330 8.605 144.630 8.625 ;
        RECT 145.300 8.605 145.600 8.625 ;
        RECT 146.250 8.605 146.550 8.615 ;
        RECT 147.220 8.605 147.520 8.625 ;
        RECT 148.170 8.605 148.470 8.625 ;
        RECT 149.130 8.605 149.430 8.625 ;
        RECT 150.100 8.605 150.400 8.625 ;
        RECT 151.050 8.605 151.350 8.625 ;
        RECT 152.030 8.605 152.330 8.635 ;
        RECT 152.980 8.605 153.280 8.625 ;
        RECT 141.580 8.265 153.540 8.605 ;
        RECT 156.390 8.515 157.330 9.365 ;
        RECT 156.410 8.490 157.310 8.515 ;
        RECT 141.580 8.235 141.920 8.265 ;
        RECT 143.370 8.235 143.670 8.265 ;
        RECT 144.330 8.235 144.630 8.265 ;
        RECT 145.300 8.235 145.600 8.265 ;
        RECT 146.250 8.225 146.550 8.265 ;
        RECT 147.220 8.235 147.520 8.265 ;
        RECT 148.170 8.235 148.470 8.265 ;
        RECT 149.130 8.235 149.430 8.265 ;
        RECT 150.100 8.235 150.400 8.265 ;
        RECT 151.050 8.235 151.350 8.265 ;
        RECT 152.030 8.245 152.330 8.265 ;
        RECT 152.980 8.235 153.280 8.265 ;
        RECT 126.705 6.610 128.155 6.630 ;
        RECT 126.680 5.110 131.220 6.610 ;
        RECT 126.705 5.090 128.155 5.110 ;
      LAYER met3 ;
        RECT 38.415 16.960 39.905 16.985 ;
        RECT 123.485 16.960 124.975 16.985 ;
        RECT 38.410 15.460 58.840 16.960 ;
        RECT 123.480 15.460 128.210 16.960 ;
        RECT 38.415 15.435 39.905 15.460 ;
        RECT 123.485 15.435 124.975 15.460 ;
        RECT 134.330 8.535 135.230 9.420 ;
        RECT 156.410 8.605 157.310 9.390 ;
        RECT 134.305 7.645 135.255 8.535 ;
        RECT 156.385 7.715 157.335 8.605 ;
        RECT 156.410 7.710 157.310 7.715 ;
        RECT 134.330 7.640 135.230 7.645 ;
        RECT 123.425 6.610 124.915 6.635 ;
        RECT 123.420 5.110 128.180 6.610 ;
        RECT 123.425 5.085 124.915 5.110 ;
      LAYER met4 ;
        RECT 3.990 223.710 4.290 224.760 ;
        RECT 7.670 223.710 7.970 224.760 ;
        RECT 11.350 223.710 11.650 224.760 ;
        RECT 15.030 223.710 15.330 224.760 ;
        RECT 18.710 223.710 19.010 224.760 ;
        RECT 22.390 223.710 22.690 224.760 ;
        RECT 26.070 223.710 26.370 224.760 ;
        RECT 29.750 223.710 30.050 224.760 ;
        RECT 33.430 223.710 33.730 224.760 ;
        RECT 37.110 223.710 37.410 224.760 ;
        RECT 40.790 223.710 41.090 224.760 ;
        RECT 44.470 223.710 44.770 224.760 ;
        RECT 48.150 223.710 48.450 224.760 ;
        RECT 51.830 223.710 52.130 224.760 ;
        RECT 55.510 223.710 55.810 224.760 ;
        RECT 59.190 223.710 59.490 224.760 ;
        RECT 62.870 223.710 63.170 224.760 ;
        RECT 66.550 223.710 66.850 224.760 ;
        RECT 70.230 223.710 70.530 224.760 ;
        RECT 73.910 223.710 74.210 224.760 ;
        RECT 77.590 223.710 77.890 224.760 ;
        RECT 81.270 223.710 81.570 224.760 ;
        RECT 84.950 223.710 85.250 224.760 ;
        RECT 88.630 223.710 88.930 224.760 ;
        RECT 2.000 222.630 90.470 223.710 ;
        RECT 49.190 220.760 50.270 222.630 ;
        RECT 57.305 16.960 58.815 16.965 ;
        RECT 2.500 15.460 39.910 16.960 ;
        RECT 57.305 15.460 124.980 16.960 ;
        RECT 57.305 15.455 58.815 15.460 ;
        RECT 50.500 5.110 124.920 6.610 ;
        RECT 134.330 1.000 135.230 8.540 ;
        RECT 156.410 1.000 157.310 8.610 ;
  END
END tt_um_Saitama224_comp
END LIBRARY

