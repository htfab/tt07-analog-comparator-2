VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Saitama224_comp
  CLASS BLOCK ;
  FOREIGN tt_um_Saitama224_comp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 73.120 197.630 76.380 209.820 ;
        RECT 77.710 206.450 82.670 211.640 ;
      LAYER pwell ;
        RECT 84.510 206.520 91.470 211.620 ;
        RECT 93.200 208.830 100.160 211.500 ;
      LAYER nwell ;
        RECT 101.520 208.850 106.480 211.640 ;
        RECT 77.715 199.985 82.675 205.175 ;
        RECT 101.500 202.370 106.460 207.560 ;
        RECT 77.700 195.910 82.660 198.700 ;
      LAYER pwell ;
        RECT 84.160 195.900 91.120 198.570 ;
        RECT 93.180 195.890 100.140 200.990 ;
      LAYER nwell ;
        RECT 101.510 195.900 106.470 201.090 ;
        RECT 108.060 197.630 111.320 209.820 ;
      LAYER li1 ;
        RECT 77.890 211.290 82.490 211.460 ;
        RECT 77.890 210.980 78.060 211.290 ;
        RECT 73.780 209.640 75.720 209.660 ;
        RECT 73.300 209.470 76.200 209.640 ;
        RECT 73.300 197.980 73.470 209.470 ;
        RECT 73.780 209.440 75.720 209.470 ;
        RECT 74.100 208.960 75.400 209.130 ;
        RECT 73.870 198.705 74.040 208.745 ;
        RECT 75.460 198.705 75.630 208.745 ;
        RECT 74.100 198.320 75.400 198.490 ;
        RECT 76.030 197.980 76.200 209.470 ;
        RECT 77.860 207.110 78.080 210.980 ;
        RECT 78.690 210.780 81.690 210.950 ;
        RECT 78.460 207.525 78.630 210.565 ;
        RECT 81.750 207.525 81.920 210.565 ;
        RECT 78.690 207.140 81.690 207.310 ;
        RECT 77.890 206.800 78.060 207.110 ;
        RECT 82.320 206.800 82.490 211.290 ;
        RECT 77.890 206.630 82.490 206.800 ;
        RECT 84.690 211.270 91.290 211.440 ;
        RECT 84.690 206.870 84.860 211.270 ;
        RECT 91.120 210.960 91.290 211.270 ;
        RECT 93.380 211.150 99.980 211.320 ;
        RECT 85.490 210.760 90.490 210.930 ;
        RECT 85.260 207.550 85.430 210.590 ;
        RECT 90.550 207.550 90.720 210.590 ;
        RECT 85.490 207.210 90.490 207.380 ;
        RECT 91.090 207.180 91.320 210.960 ;
        RECT 93.380 210.840 93.550 211.150 ;
        RECT 99.810 210.840 99.980 211.150 ;
        RECT 101.700 211.290 106.300 211.460 ;
        RECT 93.350 209.490 93.570 210.840 ;
        RECT 94.180 210.640 99.180 210.810 ;
        RECT 93.950 209.860 94.120 210.470 ;
        RECT 99.240 209.860 99.410 210.470 ;
        RECT 94.180 209.520 99.180 209.690 ;
        RECT 99.780 209.490 100.020 210.840 ;
        RECT 93.380 209.180 93.550 209.490 ;
        RECT 99.810 209.180 99.980 209.490 ;
        RECT 93.380 209.010 99.980 209.180 ;
        RECT 101.700 209.200 101.870 211.290 ;
        RECT 106.130 210.980 106.300 211.290 ;
        RECT 102.500 210.780 105.500 210.950 ;
        RECT 102.270 209.925 102.440 210.565 ;
        RECT 105.560 209.925 105.730 210.565 ;
        RECT 102.500 209.540 105.500 209.710 ;
        RECT 106.100 209.510 106.330 210.980 ;
        RECT 108.720 209.640 110.660 209.660 ;
        RECT 106.130 209.200 106.300 209.510 ;
        RECT 101.700 209.030 106.300 209.200 ;
        RECT 108.240 209.470 111.140 209.640 ;
        RECT 101.680 207.210 106.280 207.380 ;
        RECT 91.120 206.870 91.290 207.180 ;
        RECT 101.680 206.900 101.850 207.210 ;
        RECT 106.110 206.900 106.280 207.210 ;
        RECT 84.690 206.700 91.290 206.870 ;
        RECT 77.895 204.825 82.495 204.995 ;
        RECT 77.895 204.520 78.065 204.825 ;
        RECT 82.325 204.520 82.495 204.825 ;
        RECT 77.870 200.640 78.090 204.520 ;
        RECT 78.695 204.315 81.695 204.485 ;
        RECT 78.465 201.060 78.635 204.100 ;
        RECT 81.755 201.060 81.925 204.100 ;
        RECT 78.695 200.675 81.695 200.845 ;
        RECT 82.310 200.640 82.520 204.520 ;
        RECT 101.650 203.030 101.880 206.900 ;
        RECT 102.480 206.700 105.480 206.870 ;
        RECT 102.250 203.445 102.420 206.485 ;
        RECT 105.540 203.445 105.710 206.485 ;
        RECT 102.480 203.060 105.480 203.230 ;
        RECT 106.080 203.030 106.310 206.900 ;
        RECT 101.680 202.720 101.850 203.030 ;
        RECT 106.110 202.720 106.280 203.030 ;
        RECT 101.680 202.550 106.280 202.720 ;
        RECT 93.360 200.640 99.960 200.810 ;
        RECT 77.895 200.335 78.065 200.640 ;
        RECT 82.325 200.335 82.495 200.640 ;
        RECT 77.895 200.165 82.495 200.335 ;
        RECT 93.360 200.330 93.530 200.640 ;
        RECT 77.880 198.350 82.480 198.520 ;
        RECT 77.880 198.040 78.050 198.350 ;
        RECT 82.310 198.040 82.480 198.350 ;
        RECT 84.340 198.220 90.940 198.390 ;
        RECT 73.300 197.810 76.200 197.980 ;
        RECT 77.860 196.570 78.080 198.040 ;
        RECT 78.680 197.840 81.680 198.010 ;
        RECT 78.450 196.985 78.620 197.625 ;
        RECT 81.740 196.985 81.910 197.625 ;
        RECT 78.680 196.600 81.680 196.770 ;
        RECT 82.290 196.570 82.510 198.040 ;
        RECT 84.340 197.910 84.510 198.220 ;
        RECT 90.770 197.910 90.940 198.220 ;
        RECT 77.880 196.260 78.050 196.570 ;
        RECT 82.310 196.260 82.480 196.570 ;
        RECT 84.290 196.560 84.550 197.910 ;
        RECT 85.140 197.710 90.140 197.880 ;
        RECT 84.910 196.930 85.080 197.540 ;
        RECT 90.200 196.930 90.370 197.540 ;
        RECT 85.140 196.590 90.140 196.760 ;
        RECT 90.740 196.560 90.980 197.910 ;
        RECT 77.880 196.090 82.480 196.260 ;
        RECT 84.340 196.250 84.510 196.560 ;
        RECT 90.770 196.250 90.940 196.560 ;
        RECT 93.340 196.550 93.560 200.330 ;
        RECT 94.160 200.130 99.160 200.300 ;
        RECT 93.930 196.920 94.100 199.960 ;
        RECT 99.220 196.920 99.390 199.960 ;
        RECT 94.160 196.580 99.160 196.750 ;
        RECT 84.340 196.080 90.940 196.250 ;
        RECT 93.360 196.240 93.530 196.550 ;
        RECT 99.790 196.240 99.960 200.640 ;
        RECT 101.690 200.740 106.290 200.910 ;
        RECT 101.690 200.430 101.860 200.740 ;
        RECT 106.120 200.430 106.290 200.740 ;
        RECT 101.660 196.560 101.890 200.430 ;
        RECT 102.490 200.230 105.490 200.400 ;
        RECT 102.260 196.975 102.430 200.015 ;
        RECT 105.550 196.975 105.720 200.015 ;
        RECT 102.490 196.590 105.490 196.760 ;
        RECT 106.100 196.560 106.310 200.430 ;
        RECT 108.240 197.980 108.410 209.470 ;
        RECT 108.720 209.450 110.660 209.470 ;
        RECT 109.040 208.960 110.340 209.130 ;
        RECT 108.810 198.705 108.980 208.745 ;
        RECT 110.400 198.705 110.570 208.745 ;
        RECT 109.040 198.320 110.340 198.490 ;
        RECT 110.970 197.980 111.140 209.470 ;
        RECT 108.240 197.810 111.140 197.980 ;
        RECT 93.360 196.070 99.960 196.240 ;
        RECT 101.690 196.250 101.860 196.560 ;
        RECT 106.120 196.250 106.290 196.560 ;
        RECT 101.690 196.080 106.290 196.250 ;
      LAYER mcon ;
        RECT 74.180 208.960 75.320 209.130 ;
        RECT 73.870 198.785 74.040 208.665 ;
        RECT 75.460 198.785 75.630 208.665 ;
        RECT 74.180 198.320 75.320 198.490 ;
        RECT 77.860 207.110 78.080 210.980 ;
        RECT 78.770 210.780 81.610 210.950 ;
        RECT 78.460 207.605 78.630 210.485 ;
        RECT 81.750 207.605 81.920 210.485 ;
        RECT 78.770 207.140 81.610 207.310 ;
        RECT 85.570 210.760 90.410 210.930 ;
        RECT 85.260 207.630 85.430 210.510 ;
        RECT 90.550 207.630 90.720 210.510 ;
        RECT 85.570 207.210 90.410 207.380 ;
        RECT 91.090 207.180 91.320 210.960 ;
        RECT 93.350 209.490 93.570 210.840 ;
        RECT 94.260 210.640 99.100 210.810 ;
        RECT 93.950 209.940 94.120 210.390 ;
        RECT 99.240 209.940 99.410 210.390 ;
        RECT 94.260 209.520 99.100 209.690 ;
        RECT 99.780 209.490 100.020 210.840 ;
        RECT 102.580 210.780 105.420 210.950 ;
        RECT 102.270 210.005 102.440 210.485 ;
        RECT 105.560 210.005 105.730 210.485 ;
        RECT 102.580 209.540 105.420 209.710 ;
        RECT 106.100 209.510 106.330 210.980 ;
        RECT 78.775 204.315 81.615 204.485 ;
        RECT 78.465 201.140 78.635 204.020 ;
        RECT 81.755 201.140 81.925 204.020 ;
        RECT 78.775 200.675 81.615 200.845 ;
        RECT 101.650 203.030 101.880 206.900 ;
        RECT 102.560 206.700 105.400 206.870 ;
        RECT 102.250 203.525 102.420 206.405 ;
        RECT 105.540 203.525 105.710 206.405 ;
        RECT 102.560 203.060 105.400 203.230 ;
        RECT 106.080 203.030 106.310 206.900 ;
        RECT 77.860 196.570 78.080 198.040 ;
        RECT 78.760 197.840 81.600 198.010 ;
        RECT 78.450 197.065 78.620 197.545 ;
        RECT 81.740 197.065 81.910 197.545 ;
        RECT 78.760 196.600 81.600 196.770 ;
        RECT 82.290 196.570 82.510 198.040 ;
        RECT 84.290 196.560 84.550 197.910 ;
        RECT 85.220 197.710 90.060 197.880 ;
        RECT 84.910 197.010 85.080 197.460 ;
        RECT 90.200 197.010 90.370 197.460 ;
        RECT 85.220 196.590 90.060 196.760 ;
        RECT 90.740 196.560 90.980 197.910 ;
        RECT 93.340 196.550 93.560 200.330 ;
        RECT 94.240 200.130 99.080 200.300 ;
        RECT 93.930 197.000 94.100 199.880 ;
        RECT 99.220 197.000 99.390 199.880 ;
        RECT 94.240 196.580 99.080 196.750 ;
        RECT 101.660 196.560 101.890 200.430 ;
        RECT 102.570 200.230 105.410 200.400 ;
        RECT 102.260 197.055 102.430 199.935 ;
        RECT 105.550 197.055 105.720 199.935 ;
        RECT 102.570 196.590 105.410 196.760 ;
        RECT 106.100 196.560 106.310 200.430 ;
        RECT 109.120 208.960 110.260 209.130 ;
        RECT 108.810 198.785 108.980 208.665 ;
        RECT 110.400 198.785 110.570 208.665 ;
        RECT 109.120 198.320 110.260 198.490 ;
      LAYER met1 ;
        RECT 71.865 213.835 117.645 214.205 ;
        RECT 71.865 211.725 72.235 213.835 ;
        RECT 73.040 212.800 106.580 213.260 ;
        RECT 71.865 211.355 73.735 211.725 ;
        RECT 77.860 211.520 78.100 212.800 ;
        RECT 99.310 211.980 102.370 212.170 ;
        RECT 73.365 209.750 73.735 211.355 ;
        RECT 73.240 209.370 76.290 209.750 ;
        RECT 77.800 209.170 78.150 211.520 ;
        RECT 78.710 210.750 81.670 210.980 ;
        RECT 85.510 210.730 90.470 210.960 ;
        RECT 78.430 209.170 78.660 210.545 ;
        RECT 74.120 209.140 75.380 209.160 ;
        RECT 73.860 208.930 75.380 209.140 ;
        RECT 77.800 208.940 78.660 209.170 ;
        RECT 73.860 208.725 74.160 208.930 ;
        RECT 73.840 208.700 74.160 208.725 ;
        RECT 73.840 198.880 74.070 208.700 ;
        RECT 73.770 198.725 74.070 198.880 ;
        RECT 75.430 199.350 75.660 208.725 ;
        RECT 77.800 202.670 78.150 208.940 ;
        RECT 78.430 207.545 78.660 208.940 ;
        RECT 81.720 209.230 81.950 210.545 ;
        RECT 85.230 209.230 85.460 210.570 ;
        RECT 81.720 208.970 85.460 209.230 ;
        RECT 81.720 207.545 81.950 208.970 ;
        RECT 85.230 207.790 85.460 208.970 ;
        RECT 90.520 210.260 90.750 210.570 ;
        RECT 91.050 210.260 91.400 211.540 ;
        RECT 93.290 210.260 93.640 211.400 ;
        RECT 94.200 210.610 99.160 210.840 ;
        RECT 99.310 210.450 99.530 211.980 ;
        RECT 93.920 210.260 94.150 210.450 ;
        RECT 90.520 209.950 94.150 210.260 ;
        RECT 85.230 207.570 85.660 207.790 ;
        RECT 90.520 207.570 90.750 209.950 ;
        RECT 85.320 207.410 85.660 207.570 ;
        RECT 78.710 207.110 81.670 207.340 ;
        RECT 85.320 207.190 90.470 207.410 ;
        RECT 85.510 207.180 90.470 207.190 ;
        RECT 79.980 204.515 80.280 207.110 ;
        RECT 89.940 205.990 90.280 207.180 ;
        RECT 91.050 206.640 91.400 209.950 ;
        RECT 93.290 208.940 93.640 209.950 ;
        RECT 93.920 209.880 94.150 209.950 ;
        RECT 99.210 210.360 99.530 210.450 ;
        RECT 99.210 209.880 99.440 210.360 ;
        RECT 94.380 209.720 94.740 209.750 ;
        RECT 94.200 209.490 99.160 209.720 ;
        RECT 94.380 205.990 94.740 209.490 ;
        RECT 99.720 208.930 100.100 211.410 ;
        RECT 102.150 210.545 102.370 211.980 ;
        RECT 106.130 211.540 106.370 212.800 ;
        RECT 102.520 210.750 105.480 210.980 ;
        RECT 102.150 210.360 102.470 210.545 ;
        RECT 102.240 209.945 102.470 210.360 ;
        RECT 105.530 210.310 105.760 210.545 ;
        RECT 106.040 210.310 106.410 211.540 ;
        RECT 105.530 210.100 106.410 210.310 ;
        RECT 105.530 209.945 105.760 210.100 ;
        RECT 102.520 209.510 105.480 209.740 ;
        RECT 89.940 205.620 94.740 205.990 ;
        RECT 89.940 205.610 90.280 205.620 ;
        RECT 78.715 204.500 81.675 204.515 ;
        RECT 78.715 204.285 81.940 204.500 ;
        RECT 81.610 204.080 81.940 204.285 ;
        RECT 78.435 202.670 78.665 204.080 ;
        RECT 81.610 203.840 81.955 204.080 ;
        RECT 77.800 202.450 78.665 202.670 ;
        RECT 77.800 200.110 78.150 202.450 ;
        RECT 78.435 201.080 78.665 202.450 ;
        RECT 81.725 201.080 81.955 203.840 ;
        RECT 78.715 200.645 81.675 200.875 ;
        RECT 79.980 199.350 80.280 200.645 ;
        RECT 75.430 199.090 80.280 199.350 ;
        RECT 75.430 198.725 75.660 199.090 ;
        RECT 73.770 194.830 73.970 198.725 ;
        RECT 74.120 198.290 75.380 198.520 ;
        RECT 77.800 197.410 78.150 198.570 ;
        RECT 79.980 198.040 80.280 199.090 ;
        RECT 78.700 197.810 81.660 198.040 ;
        RECT 78.420 197.410 78.650 197.605 ;
        RECT 77.800 197.200 78.650 197.410 ;
        RECT 77.800 196.050 78.150 197.200 ;
        RECT 78.420 197.005 78.650 197.200 ;
        RECT 81.710 197.310 81.940 197.605 ;
        RECT 81.710 197.005 82.050 197.310 ;
        RECT 78.700 196.570 81.660 196.800 ;
        RECT 81.810 195.740 82.050 197.005 ;
        RECT 82.250 196.000 82.570 205.110 ;
        RECT 99.770 203.920 100.040 208.930 ;
        RECT 84.260 203.580 100.040 203.920 ;
        RECT 84.260 198.470 84.580 203.580 ;
        RECT 89.880 201.540 94.680 201.910 ;
        RECT 84.210 196.010 84.600 198.470 ;
        RECT 89.880 197.910 90.240 201.540 ;
        RECT 85.160 197.780 90.240 197.910 ;
        RECT 85.160 197.680 90.120 197.780 ;
        RECT 84.880 197.310 85.110 197.520 ;
        RECT 84.760 196.950 85.110 197.310 ;
        RECT 90.170 197.420 90.400 197.520 ;
        RECT 90.700 197.420 91.070 198.470 ;
        RECT 93.280 197.420 93.600 200.920 ;
        RECT 94.340 200.330 94.680 201.540 ;
        RECT 94.180 200.320 99.140 200.330 ;
        RECT 94.180 200.100 99.380 200.320 ;
        RECT 99.040 199.940 99.380 200.100 ;
        RECT 93.900 197.420 94.130 199.940 ;
        RECT 99.040 199.830 99.420 199.940 ;
        RECT 90.170 197.110 94.130 197.420 ;
        RECT 90.170 196.950 90.400 197.110 ;
        RECT 84.760 195.740 85.000 196.950 ;
        RECT 85.160 196.560 90.120 196.790 ;
        RECT 90.700 196.000 91.070 197.110 ;
        RECT 81.810 195.480 85.000 195.740 ;
        RECT 83.570 195.090 83.990 195.480 ;
        RECT 91.800 194.830 92.260 197.110 ;
        RECT 93.280 196.010 93.600 197.110 ;
        RECT 93.900 196.940 94.130 197.110 ;
        RECT 99.190 197.190 99.420 199.830 ;
        RECT 99.190 196.940 99.600 197.190 ;
        RECT 94.180 196.550 99.140 196.780 ;
        RECT 99.380 195.720 99.600 196.940 ;
        RECT 101.600 196.000 101.960 207.480 ;
        RECT 103.690 206.900 103.990 209.510 ;
        RECT 102.500 206.670 105.460 206.900 ;
        RECT 102.220 203.740 102.450 206.465 ;
        RECT 105.510 205.040 105.740 206.465 ;
        RECT 106.040 205.040 106.410 210.100 ;
        RECT 110.660 211.030 117.540 211.390 ;
        RECT 110.660 209.710 111.020 211.030 ;
        RECT 108.160 209.350 111.210 209.710 ;
        RECT 109.060 209.110 110.320 209.160 ;
        RECT 109.060 208.930 110.590 209.110 ;
        RECT 110.290 208.725 110.590 208.930 ;
        RECT 105.510 204.840 106.410 205.040 ;
        RECT 102.220 203.465 102.590 203.740 ;
        RECT 105.510 203.465 105.740 204.840 ;
        RECT 102.260 203.260 102.590 203.465 ;
        RECT 102.260 203.080 105.460 203.260 ;
        RECT 102.500 203.030 105.460 203.080 ;
        RECT 104.040 201.760 104.340 203.030 ;
        RECT 106.040 202.460 106.410 204.840 ;
        RECT 108.780 201.760 109.010 208.725 ;
        RECT 110.290 208.670 110.600 208.725 ;
        RECT 104.040 201.500 109.010 201.760 ;
        RECT 104.040 200.430 104.340 201.500 ;
        RECT 102.510 200.200 105.470 200.430 ;
        RECT 102.230 197.190 102.460 199.995 ;
        RECT 102.140 196.995 102.460 197.190 ;
        RECT 105.520 198.590 105.750 199.995 ;
        RECT 106.050 198.590 106.390 200.990 ;
        RECT 108.780 198.725 109.010 201.500 ;
        RECT 110.370 198.890 110.600 208.670 ;
        RECT 110.370 198.725 110.690 198.890 ;
        RECT 105.520 198.390 106.390 198.590 ;
        RECT 105.520 196.995 105.750 198.390 ;
        RECT 102.140 195.720 102.360 196.995 ;
        RECT 102.510 196.560 105.470 196.790 ;
        RECT 106.050 195.990 106.390 198.390 ;
        RECT 109.060 198.290 110.320 198.520 ;
        RECT 99.380 195.460 102.360 195.720 ;
        RECT 110.490 194.830 110.690 198.725 ;
        RECT 73.160 194.300 111.310 194.830 ;
      LAYER via ;
        RECT 117.350 213.890 117.610 214.150 ;
        RECT 73.260 212.800 73.720 213.260 ;
        RECT 83.640 195.150 83.910 195.410 ;
        RECT 117.150 211.060 117.420 211.350 ;
        RECT 75.000 194.390 75.370 194.720 ;
      LAYER met2 ;
        RECT 117.240 213.810 117.700 214.230 ;
        RECT 40.725 212.610 73.870 213.480 ;
        RECT 117.030 210.980 117.540 211.420 ;
        RECT 83.520 195.050 84.090 195.540 ;
        RECT 74.790 194.170 75.580 194.940 ;
      LAYER via2 ;
        RECT 117.300 213.880 117.610 214.170 ;
        RECT 41.250 212.780 41.850 213.330 ;
        RECT 117.130 211.050 117.440 211.370 ;
        RECT 83.620 195.140 83.930 195.430 ;
        RECT 74.880 194.300 75.480 194.830 ;
      LAYER met3 ;
        RECT 117.200 213.780 117.760 214.310 ;
        RECT 40.700 212.480 42.290 213.580 ;
        RECT 117.110 211.030 117.460 211.390 ;
        RECT 83.490 195.030 84.120 195.560 ;
        RECT 74.700 194.070 75.680 195.020 ;
      LAYER via3 ;
        RECT 117.260 213.860 117.630 214.190 ;
        RECT 41.190 212.730 41.910 213.360 ;
        RECT 83.600 195.120 83.950 195.450 ;
        RECT 74.850 194.230 75.520 194.870 ;
      LAYER met4 ;
        RECT 4.290 224.870 7.670 225.460 ;
        RECT 7.970 224.870 11.350 225.460 ;
        RECT 11.650 224.870 15.030 225.460 ;
        RECT 15.330 224.870 18.710 225.460 ;
        RECT 19.010 224.870 22.390 225.460 ;
        RECT 22.690 224.870 26.070 225.460 ;
        RECT 26.370 224.870 29.750 225.460 ;
        RECT 30.050 224.870 33.430 225.460 ;
        RECT 33.730 224.870 37.110 225.460 ;
        RECT 37.410 224.870 40.790 225.460 ;
        RECT 41.090 224.870 44.470 225.460 ;
        RECT 44.770 224.870 48.150 225.460 ;
        RECT 48.450 224.870 51.830 225.460 ;
        RECT 52.130 224.870 55.510 225.460 ;
        RECT 55.810 224.870 59.190 225.460 ;
        RECT 59.490 224.870 62.870 225.460 ;
        RECT 62.665 224.760 62.870 224.870 ;
        RECT 63.170 224.870 66.550 225.460 ;
        RECT 66.850 224.870 70.230 225.460 ;
        RECT 70.530 224.870 73.910 225.460 ;
        RECT 74.210 224.870 77.590 225.460 ;
        RECT 77.890 224.870 81.270 225.460 ;
        RECT 81.570 224.870 84.950 225.460 ;
        RECT 85.250 224.870 88.630 225.460 ;
        RECT 63.170 224.760 63.255 224.870 ;
        RECT 2.500 212.350 42.470 213.850 ;
        RECT 62.665 195.250 63.255 224.760 ;
        RECT 84.950 224.750 85.250 224.760 ;
        RECT 88.630 224.750 88.930 224.760 ;
        RECT 147.510 224.740 147.810 224.760 ;
        RECT 116.740 213.580 157.310 214.480 ;
        RECT 116.900 210.760 135.230 211.660 ;
        RECT 50.500 193.750 75.990 195.250 ;
        RECT 83.390 191.500 84.230 195.640 ;
        RECT 83.390 190.600 113.150 191.500 ;
        RECT 112.250 1.000 113.150 190.600 ;
        RECT 134.330 1.000 135.230 210.760 ;
        RECT 156.410 1.000 157.310 213.580 ;
  END
END tt_um_Saitama224_comp
END LIBRARY

