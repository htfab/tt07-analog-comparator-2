magic
tech sky130A
magscale 1 2
timestamp 1716851390
<< pwell >>
rect 17064 41438 17132 41558
rect 19808 39966 19876 40064
<< locali >>
rect 14756 41888 15144 41932
rect 21744 41890 22132 41932
<< viali >>
rect 15572 41422 15616 42196
rect 18218 41436 18264 42192
rect 18670 41898 18714 42168
rect 19956 41898 20004 42168
rect 21220 41902 21266 42196
rect 15574 40128 15618 40904
rect 16462 40128 16504 40904
rect 20330 40606 20376 41380
rect 21216 40606 21262 41380
rect 15572 39314 15616 39608
rect 16458 39314 16502 39608
rect 16858 39312 16910 39582
rect 18148 39312 18196 39582
rect 18668 39310 18712 40066
rect 20332 39312 20378 40086
rect 21220 39312 21262 40086
<< metal1 >>
rect 14373 42830 23529 42841
rect 14373 42778 23470 42830
rect 23522 42778 23529 42830
rect 14373 42767 23529 42778
rect 14373 42345 14447 42767
rect 14608 42560 14652 42652
rect 14744 42560 21316 42652
rect 14373 42271 14747 42345
rect 15572 42304 15620 42560
rect 19862 42396 20474 42434
rect 14673 41950 14747 42271
rect 15560 42196 15630 42304
rect 14648 41874 15258 41950
rect 14772 41740 14832 41828
rect 15560 41422 15572 42196
rect 15616 41834 15630 42196
rect 18210 42192 18280 42308
rect 18210 42052 18218 42192
rect 18130 41990 18218 42052
rect 15616 41788 15722 41834
rect 16366 41794 17070 41846
rect 15616 41422 15630 41788
rect 15560 40904 15630 41422
rect 15560 40128 15574 40904
rect 15618 40534 15630 40904
rect 15996 40882 16056 41458
rect 17064 41438 17132 41558
rect 17988 41198 18056 41466
rect 18210 41436 18218 41990
rect 18264 42052 18280 42192
rect 18658 42168 18728 42280
rect 18658 42052 18670 42168
rect 18264 41990 18670 42052
rect 18264 41436 18280 41990
rect 18658 41898 18670 41990
rect 18714 42052 18728 42168
rect 19862 42072 19906 42396
rect 19944 42168 20020 42282
rect 18714 41990 18802 42052
rect 18714 41898 18728 41990
rect 18658 41788 18728 41898
rect 18210 41328 18280 41436
rect 18876 41198 18948 41950
rect 19944 41898 19956 42168
rect 20004 41898 20020 42168
rect 20430 42072 20474 42396
rect 21226 42308 21274 42560
rect 21208 42196 21282 42308
rect 21208 42062 21220 42196
rect 21120 42020 21220 42062
rect 19944 41786 20020 41898
rect 17988 41124 18948 41198
rect 17988 41122 18056 41124
rect 16450 40904 16514 41022
rect 16322 40768 16388 40900
rect 15618 40490 15718 40534
rect 15618 40128 15630 40490
rect 15560 40022 15630 40128
rect 15996 39870 16056 40152
rect 15110 39818 16056 39870
rect 14754 38966 14794 39776
rect 15560 39608 15630 39714
rect 15560 39314 15572 39608
rect 15616 39482 15630 39608
rect 15996 39576 16056 39818
rect 16450 40128 16462 40904
rect 16504 40128 16514 40904
rect 19954 40784 20008 41786
rect 16450 39608 16514 40128
rect 16852 40716 20008 40784
rect 20320 41380 20392 41496
rect 16852 39694 16916 40716
rect 20320 40606 20330 41380
rect 20376 40606 20392 41380
rect 20738 41362 20798 41938
rect 21208 41902 21220 42020
rect 21266 41902 21282 42196
rect 22132 42270 23508 42278
rect 22132 42212 23430 42270
rect 23484 42212 23508 42270
rect 22132 42206 23508 42212
rect 22132 41942 22204 42206
rect 21208 41380 21282 41902
rect 21632 41870 22242 41942
rect 22058 41734 22118 41822
rect 21208 41008 21216 41380
rect 21116 40968 21216 41008
rect 20452 40616 20518 40748
rect 17976 40308 18936 40382
rect 15616 39440 15712 39482
rect 15616 39314 15630 39440
rect 15560 39210 15630 39314
rect 16362 39148 16410 39462
rect 16450 39314 16458 39608
rect 16502 39314 16514 39608
rect 16450 39200 16514 39314
rect 16842 39582 16920 39694
rect 16842 39312 16858 39582
rect 16910 39312 16920 39582
rect 17976 39556 18048 40308
rect 18656 40066 18720 40184
rect 18140 39582 18214 39694
rect 18140 39484 18148 39582
rect 16842 39202 16920 39312
rect 16952 39148 17000 39462
rect 18058 39422 18148 39484
rect 18140 39312 18148 39422
rect 18196 39484 18214 39582
rect 18656 39484 18668 40066
rect 18196 39422 18668 39484
rect 18196 39312 18214 39422
rect 18140 39200 18214 39312
rect 16362 39096 17000 39148
rect 16714 39082 16798 39096
rect 16714 39030 16728 39082
rect 16782 39030 16798 39082
rect 16714 39018 16798 39030
rect 18360 38966 18452 39422
rect 18656 39310 18668 39422
rect 18712 39484 18720 40066
rect 18868 40038 18936 40308
rect 20320 40086 20392 40606
rect 19808 39966 19876 40064
rect 18712 39422 18806 39484
rect 18712 39310 18720 39422
rect 18656 39202 18720 39310
rect 19876 39144 19920 39438
rect 20320 39312 20332 40086
rect 20378 39312 20392 40086
rect 20808 40352 20868 40638
rect 21208 40606 21216 40968
rect 21262 40606 21282 41380
rect 21208 40492 21282 40606
rect 20808 40300 21786 40352
rect 20808 40062 20868 40300
rect 21210 40086 21278 40198
rect 21210 39718 21220 40086
rect 21118 39678 21220 39718
rect 20320 39200 20392 39312
rect 20428 39144 20472 39438
rect 21210 39312 21220 39678
rect 21262 39312 21278 40086
rect 21210 39198 21278 39312
rect 19876 39092 20472 39144
rect 22098 38966 22138 39778
rect 14632 38944 22262 38966
rect 14632 38878 15000 38944
rect 15074 38878 22262 38944
rect 14632 38860 22262 38878
<< via1 >>
rect 23470 42778 23522 42830
rect 14652 42560 14744 42652
rect 23430 42212 23484 42270
rect 16728 39030 16782 39082
rect 15000 38878 15074 38944
<< metal2 >>
rect 23448 42834 23540 42846
rect 23448 42776 23460 42834
rect 23522 42776 23540 42834
rect 23448 42762 23540 42776
rect 8145 42666 14774 42696
rect 8145 42556 8250 42666
rect 8370 42652 14774 42666
rect 8370 42560 14652 42652
rect 14744 42560 14774 42652
rect 8370 42556 14774 42560
rect 8145 42522 14774 42556
rect 23406 42274 23508 42284
rect 23406 42210 23426 42274
rect 23488 42210 23508 42274
rect 23406 42196 23508 42210
rect 16704 39086 16818 39108
rect 16704 39028 16724 39086
rect 16786 39028 16818 39086
rect 16704 39010 16818 39028
rect 14958 38966 15116 38988
rect 14958 38860 14976 38966
rect 15096 38860 15116 38966
rect 14958 38834 15116 38860
<< via2 >>
rect 23460 42830 23522 42834
rect 23460 42778 23470 42830
rect 23470 42778 23522 42830
rect 23460 42776 23522 42778
rect 8250 42556 8370 42666
rect 23426 42270 23488 42274
rect 23426 42212 23430 42270
rect 23430 42212 23484 42270
rect 23484 42212 23488 42270
rect 23426 42210 23488 42212
rect 16724 39082 16786 39086
rect 16724 39030 16728 39082
rect 16728 39030 16782 39082
rect 16782 39030 16786 39082
rect 16724 39028 16786 39030
rect 14976 38944 15096 38966
rect 14976 38878 15000 38944
rect 15000 38878 15074 38944
rect 15074 38878 15096 38944
rect 14976 38860 15096 38878
<< metal3 >>
rect 23440 42838 23552 42862
rect 23440 42772 23452 42838
rect 23526 42772 23552 42838
rect 23440 42756 23552 42772
rect 8140 42672 8458 42716
rect 8140 42546 8238 42672
rect 8382 42546 8458 42672
rect 8140 42496 8458 42546
rect 16698 39090 16824 39112
rect 16698 39024 16720 39090
rect 16790 39024 16824 39090
rect 16698 39006 16824 39024
rect 14940 38974 15136 39004
rect 14940 38846 14970 38974
rect 15104 38846 15136 38974
rect 14940 38814 15136 38846
<< rmetal3 >>
rect 23400 42278 23514 42290
rect 23400 42206 23422 42278
rect 23492 42206 23514 42278
rect 23400 42190 23514 42206
<< via3 >>
rect 23452 42834 23526 42838
rect 23452 42776 23460 42834
rect 23460 42776 23522 42834
rect 23522 42776 23526 42834
rect 23452 42772 23526 42776
rect 8238 42666 8382 42672
rect 8238 42556 8250 42666
rect 8250 42556 8370 42666
rect 8370 42556 8382 42666
rect 8238 42546 8382 42556
rect 23422 42274 23492 42278
rect 23422 42210 23426 42274
rect 23426 42210 23488 42274
rect 23488 42210 23492 42274
rect 23422 42206 23492 42210
rect 16720 39086 16790 39090
rect 16720 39028 16724 39086
rect 16724 39028 16786 39086
rect 16786 39028 16790 39086
rect 16720 39024 16790 39028
rect 14970 38966 15104 38974
rect 14970 38860 14976 38966
rect 14976 38860 15096 38966
rect 15096 38860 15104 38966
rect 14970 38846 15104 38860
<< metal4 >>
rect 798 45092 858 45152
rect 1534 45092 1594 45152
rect 2270 45092 2330 45152
rect 3006 45092 3066 45152
rect 3742 45092 3802 45152
rect 4478 45092 4538 45152
rect 5214 45092 5274 45152
rect 5950 45092 6010 45152
rect 6686 45092 6746 45152
rect 7422 45092 7482 45152
rect 8158 45092 8218 45152
rect 8894 45092 8954 45152
rect 9630 45092 9690 45152
rect 10366 45092 10426 45152
rect 11102 45092 11162 45152
rect 11838 45092 11898 45152
rect 12574 45092 12634 45152
rect 13310 45092 13370 45152
rect 14046 45092 14106 45152
rect 14782 45092 14842 45152
rect 15518 45092 15578 45152
rect 16254 45092 16314 45152
rect 16990 45092 17050 45152
rect 17726 45092 17786 45152
rect 798 44974 17786 45092
rect 798 44952 858 44974
rect 1534 44952 1594 44974
rect 2270 44952 2330 44974
rect 3006 44952 3066 44974
rect 3742 44952 3802 44974
rect 4478 44952 4538 44974
rect 5214 44952 5274 44974
rect 5950 44952 6010 44974
rect 6686 44952 6746 44974
rect 7422 44952 7482 44974
rect 8158 44952 8218 44974
rect 8894 44952 8954 44974
rect 9630 44952 9690 44974
rect 10366 44952 10426 44974
rect 11102 44952 11162 44974
rect 11838 44952 11898 44974
rect 200 42770 500 44152
rect 200 42672 8494 42770
rect 200 42546 8238 42672
rect 8382 42546 8494 42672
rect 200 42470 8494 42546
rect 200 1000 500 42470
rect 9800 39050 10100 44152
rect 12533 39050 12651 44974
rect 13310 44952 13370 44974
rect 14046 44952 14106 44974
rect 14782 44952 14842 44974
rect 15518 44952 15578 44974
rect 16254 44952 16314 44974
rect 16990 44950 17050 44974
rect 17726 44950 17786 44974
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44948 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 23348 42838 31462 42896
rect 23348 42772 23452 42838
rect 23526 42772 31462 42838
rect 23348 42716 31462 42772
rect 23380 42278 27046 42332
rect 23380 42206 23422 42278
rect 23492 42206 27046 42278
rect 23380 42152 27046 42206
rect 16678 39090 16846 39128
rect 9800 38974 15198 39050
rect 9800 38846 14970 38974
rect 15104 38846 15198 38974
rect 9800 38750 15198 38846
rect 16678 39024 16720 39090
rect 16790 39024 16846 39090
rect 9800 1000 10100 38750
rect 16678 38300 16846 39024
rect 16678 38120 22630 38300
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 38120
rect 26866 0 27046 42152
rect 31282 0 31462 42716
use sky130_fd_pr__nfet_01v8_HXU4AK  sky130_fd_pr__nfet_01v8_HXU4AK_0 ~/Desktop/MNEL
timestamp 1713891343
transform 1 0 19336 0 1 42033
box -696 -267 696 267
use sky130_fd_pr__nfet_01v8_HXU4AK  sky130_fd_pr__nfet_01v8_HXU4AK_1
timestamp 1713891343
transform 1 0 17528 0 1 39447
box -696 -267 696 267
use sky130_fd_pr__nfet_01v8_MXF53G  sky130_fd_pr__nfet_01v8_MXF53G_0 ~/Desktop/MNEL
timestamp 1713891343
transform 1 0 19332 0 1 39688
box -696 -510 696 510
use sky130_fd_pr__nfet_01v8_MXF53G  sky130_fd_pr__nfet_01v8_MXF53G_1
timestamp 1713891343
transform 1 0 17598 0 1 41814
box -696 -510 696 510
use sky130_fd_pr__pfet_01v8_GE7BQD  sky130_fd_pr__pfet_01v8_GE7BQD_0 ~/Desktop/MNEL
timestamp 1713898952
transform 1 0 14950 0 1 40745
box -326 -1219 326 1219
use sky130_fd_pr__pfet_01v8_GE7BQD  sky130_fd_pr__pfet_01v8_GE7BQD_1
timestamp 1713898952
transform 1 0 21938 0 1 40745
box -326 -1219 326 1219
use sky130_fd_pr__pfet_01v8_KDYT8F  sky130_fd_pr__pfet_01v8_KDYT8F_0 ~/Desktop/MNEL
timestamp 1713888985
transform 1 0 20800 0 1 42049
box -496 -279 496 279
use sky130_fd_pr__pfet_01v8_KDYT8F  sky130_fd_pr__pfet_01v8_KDYT8F_1
timestamp 1713888985
transform 1 0 16036 0 1 39461
box -496 -279 496 279
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_0 ~/Desktop/MNEL
timestamp 1713888985
transform -1 0 16039 0 -1 40516
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_1
timestamp 1713888985
transform -1 0 20798 0 -1 39699
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_2
timestamp 1713888985
transform -1 0 16038 0 -1 41809
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_3
timestamp 1713888985
transform -1 0 20796 0 -1 40993
box -496 -519 496 519
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
